interface arb_if(input clk);
   logic reset;
   logic [1:0] grant,request;
endinterface

